// ADD HAZARD DETECTION UNIT HERE!!!!

module decode (
    input clk,
    input rst_n,
    
    // Inputs from Fetch/Decode pipeline register
    input [32:0] D_in,
    
    // branch resolution signals to go back to F stage
    output flush,
    output stall,
    output [15:0] branch_target

    // pipeline data and control signals
    output [86:0] D_out;

);
    
    // internal signals from Fetch
    wire [15:0] FD_pc_plus_2;
    wire [15:0] FD_instruction;

    // declare all wire connections for decode stage
    wire [3:0] rr1_reg;               // Read register 1 selector
    wire [3:0] rr2_reg;               // Read register 2 selector
    wire [3:0] wr_reg;                // Write register selector
    wire [15:0] rr1_data;             // Data from rs register
    wire [15:0] rr2_data;             // Data from rt register
    wire [15:0] imm_value;            // Immediate value for ALU
    wire [15:0] write_data;           // Data to write to rd register

    // control signals from control module
    wire RR1Mux;                      // Read register 1 mux control
    wire RR2Mux;                      // Read register 2 mux control
    wire [1:0] ImmMux;                // Immediate value mux control
    wire ALUSrcMux;                   // ALU source mux control
    wire MemtoRegMux;                 // Memory to register mux control
    wire PCSMux;                      // PC save mux control
    wire HaltMux;                     // Halt mux control
    wire BranchRegMux;                // Branch register mux control
    wire BranchMux;                   // Branch immediate mux control
    wire RegWrite;                    // Register write control
    wire MemWrite;                    // Memory write control
    wire MemRead;                     // Enable using data memory
    wire Flag_Enable;                 // enables FF for flags
    wire ALUop;                       // bits [15:12] of inst for alu operation


    // break up the FD pipeline data
    assign FD_pc_plus_2 = D_in[31:16];    // PC + 2 forwarded to D stage
    assign FD_instruction = D_in[15:0];   // Instruction forwarded to D stage
 
    // Control unit instantiation
    control ctrl_unit(
        .instruction(FD_instruction),
        .RR1Mux(RR1Mux),
        .RR2Mux(RR2Mux),
        .ImmMux(ImmMux),
        .ALUSrcMux(ALUSrcMux),
        .MemtoRegMux(MemtoRegMux),
        .PCSMux(PCSMux),
        .HaltMux(HaltMux),
        .BranchRegMux(BranchRegMux),
        .BranchMux(BranchMux),
        .RegWrite(RegWrite),
        .MemWrite(MemWrite),
        .MemRead(MemRead),
        .Flag_Enable(Flag_Enable),
        .ALUop(ALUop)
    );

    // Register selection logic
    assign rr1_reg = RR1Mux ? FD_instruction[11:8] : FD_instruction[7:4];    // 1 : LLB / LHB , 0 : else
    assign rr2_reg = (MemWrite | MemRead) ? FD_instruction[11:8] : FD_instruction[3:0]; // LW and SW
    assign wr_reg = FD_instruction[11:8]; 

    // assign write data, data out from from writeback stage
    assign write_data = PCSMux ? FD_pc_plus_2 : data_out;
    
    // RegisterFile instantiation
    RegisterFile RF(
        .clk(clk),
        .rst(~rst_n),                  // Convert active-low to active-high
        .SrcReg1(rr1_reg),
        .SrcReg2(rr2_reg),
        .DstReg(wr_reg),
        .WriteReg(RegWrite),
        .DstData(write_data),
        .SrcData1(rr1_data),
        .SrcData2(rr2_data)
    );
    
    // Immediate value selection - based on your control logic
    assign imm_value = (ImmMux == 2'b00) ? {{12{1'b0}}, FD_instruction[3:0]} :             // 4-bit immediate (SLL, SRA, ROR)
                       (ImmMux == 2'b01) ? {{11{FD_instruction[3]}}, FD_instruction[3:0], 1'b0} : // 4-bit offset shifted (LW, SW)
                       {{8{1'b0}}, FD_instruction[7:0]};                                     // 8-bit immediate (LLB, LHB) - 2'b10
    
    // Branch resolution - using the same logic from your single-cycle implementation
    branch branch_unit(
        .branch_condition(FD_instruction[11:9]),
        .flag_reg(flags),
        .branch_taken(branch_taken)
    );
    
    // Calculate branch target
    wire [15:0] branch_value
    wire [15:0] extended_imm;
    assign extended_imm = {{6{FD_instruction[8]}}, FD_instruction[8:0], 1'b0}; // Sign-extend and shift left
    adder_16bit branch_adder(
        .A(FD_pc_plus_2),
        .B(extended_imm),
        .Sub(1'b0),
        .Sum(branch_value)
    );


    // these will actual come from hazard detection unit //
    assign stall:

    // assign flush so PC can load in the new branch addr
    assign flush = (BranchRegMux & branch_taken) | (BranchMux & branch_taken);

    // assign branch tagret, if branchMux high take output of branch_addr else take rr1 data
    assign branch_target = BranchMux ? branch_value : rr1_data;

    // assign the D_data and D_Control that goes into D/X pipe reg


    // Data signals concatenation
    wire [75:0] D_data;
    assign D_data = {
        rr1_data,     // [75:60] Data from rr1 register (16 bits)
        rr2_data,     // [59:44] Data from rr2 register (16 bits)
        write_data,   // [43:28] Data to write to wr register (16 bits)
        imm_value,    // [27:12] Immediate value from instruction (16 bits)
        rr1_reg,      // [11:8] Read register 1 number (4 bits)
        rr2_reg,      // [7:4] Read register 2 number (4 bits)
        wr_reg        // [3:0] Write register number (4 bits)
    };

    // Control signals concatenation
    wire [11:0] D_control;
    assign D_control = {
        ALUop,        // [11:8] Opcode from instruction (4 bits)
        ALUSrcMux,    // [7] ALU source selection for EX stage (1 bit)
        MemtoRegMux,  // [6] Selects memory vs. ALU result in WB (1 bit)
        PCSMux,       // [5] Selects PC+2 for PCS instructions in WB (1 bit)
        RegWrite,     // [4] Register write enable for WB (1 bit)
        MemWrite,     // [3] Memory write enable for MEM stage (1 bit)
        MemRead,      // [2] Memory read enable for MEM stage (1 bit)
        Flag_Enable,  // [1] Flag update enable for EX stage (1 bit)
        HaltMux       // [0] Halt signal (1 bit)
    };

    
    // D_out Signal Guide
    // assign final D_out with data and control values
    // 
    // [87:12] D_data (76 bits) - Data path signals
    //   [87:72] rr1_data     - Data from first source register (16 bits)
    //   [71:56] rr2_data     - Data from second source register (16 bits)
    //   [55:40] write_data   - Data to write to destination register (16 bits)
    //   [39:24] imm_value    - Immediate value from instruction (16 bits)
    //   [23:20] rr1_reg      - First source register number (4 bits)
    //   [19:16] rr2_reg      - Second source register number (4 bits)
    //   [15:12] wr_reg       - Destination register number (4 bits)
    //
    // [11:0] D_control (12 bits) - Control signals
    //   [11:8] ALUop        - ALU operation code (4 bits)
    //   [7]    ALUSrcMux    - Selects register (0) or immediate (1) for ALU B input
    //   [6]    MemtoRegMux  - Selects ALU result (0) or memory data (1) for register write
    //   [5]    PCSMux       - Selects PC+2 as write data for PCS instruction
    //   [4]    RegWrite     - Enable signal for register file writing
    //   [3]    MemWrite     - Enable signal for memory writing (SW)
    //   [2]    MemRead      - Enable signal for memory reading (LW)
    //   [1]    Flag_Enable  - Enable signal for updating ALU flags
    //   [0]    HaltMux      - Signal to halt processor execution
    
    assign D_out = {D_data, D_control}



endmodule