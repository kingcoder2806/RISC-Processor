module fetch(
    input clk,                    // Clock signal
    input rst_n,                  // Reset signal (active low)
    input stall,                  // Stall signal from hazard detection from cpu
    input flush,                  // Flush signal when branch is taken from decode
    input [15:0] branch_target,   // Branch target from ID stage
    input [15:0] cache_instruction, // From mem module in cpu
    
    // Outputs - just the basic values
    output [15:0] pc,             // Current PC value (for CPU output)
    output [31:0] F_out   // data to be passed to the FD pipe reg
);

    // Internal wires
    wire [15:0] pc_next;          // Next PC value
    wire [15:0] pc_plus_2;        // pc plus 2
    wire [15:0] instruction;
    wire halt_PC;

     // PC register logic to enable
    wire pc_en;
    assign pc_en = ~(stall);

    // PC selection logic for predict-not-taken
    // Note: Stall comes from hazard in X , flush comes from branch resolution in D, halt coms from writeback
    assign pc_next = (halt_PC & !flush)? pc :     // Halt: freeze PC unless in branch shadow!
                 flush ? branch_target :        // Branch taken: jump to target
                 pc_plus_2;                      // Normal: increment PC

    pc_reg PC(
        .clk(clk),
        .rst_n(~rst_n),
        .wen(pc_en),
        .pc_next(pc_next),
        .pc(pc)
    );

    // PC + 2 adder (for normal sequential execution)
    adder_16bit pc_incrementer(
        .A(pc),
        .B(16'h0002),
        .Sub(1'b0),
        .Sum(pc_plus_2)
    );

    // Instruction memory (removed in phase 3 since we get inst from ICache now)
    /*
    memory1c IMEM(
        .data_out(instruction),   // Output: instruction fetched
        .data_in(16'h0000),       // Not used (we don't write to instruction memory)
        .addr(pc),                // Address: current PC
        .enable(1'b1),            // Always enabled
        .wr(1'b0),                // Never write
        .clk(clk),
        .rst(~rst_n)              // Convert active-low to active-high
    );
    */

    // assign instruction from ICache inst from input
    assign instruction = cache_instruction;

    // assign halt_PC logic 
    assign halt_PC = &instruction[15:12];

    // assign data that will go into pipeline to decode
    // FD_in : {[31:16]pc_plus_2, [15:0]instruction}

    assign F_out = {pc_plus_2, instruction};

endmodule